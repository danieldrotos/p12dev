`timescale 1ns / 1ps

module mem(A, 
           CLK, 
           CS, 
           I, 
           WR, 
           CSO, 
           O);

    input [31:0] A;
    input CLK;
    input CS;
    input [31:0] I;
    input WR;
   output CSO;
   output [31:0] O;
   
   wire H;
   wire L;
   
   RAMB16_S36 #( 
      .INIT(36'h000000000), 
// //; SYMBOLS
// //; 0000c000 timer_ctrl
// //; 0000c001 timer_ar
// //; 0000c002 timer_cntr
// //; 0000c003 timer_stat
// //; 0000f000 display
// //; 0000f001 led
// //; 0000f002 portc
// //; 0000f003 portd
// //; 00000012 cyc
// //; CODE
// 0400c000 //;0000 ldl0	r0,timer_ctrl
// 0410c001 //;0001 ldl0	r1,timer_ar
// 0420c003 //;0002 ldl0	r2,timer_stat
// 0430c002 //;0003 ldl0	r3,timer_cntr
// 0440f000 //;0004 ldl0	r4,display
// 0450f001 //;0005 ldl0	r5,led
// 0460f002 //;0006 ldl0	r6,portc
// 0470f003 //;0007 ldl0	r7,portd
      .INIT_00(256'h0470f003_0460f002_0450f001_0440f000_0430c002_0420c003_0410c001_0400c000),
// 04800002 //;0008 ldl0	r8,2
// 04900000 //;0009 ldl0	r9,0		
// 02950000 //;000a st	r9,r5
// 02960000 //;000b st	r9,r6
// 02970000 //;000c st	r9,r7
// 0590a120 //;000d ldl	r9,500000	
// 06900007 //;000e ldh	r9,500000
// 02910000 //;000f st	r9,r1
      .INIT_01(256'h02910000_06900007_0590a120_02970000_02960000_02950000_04900000_04800002),
// 04a00003 //;0010 ldl0	r10,3		
// 02a00000 //;0011 st	r10,r0
// 01b60000 //;0012 ld	r11,r6
// 07bb0200 //;0013 inc	r11		
// 02b60000 //;0014 st	r11,r6		
// 01930000 //;0015 ld	r9,r3		
// 02940000 //;0016 st	r9,r4		
// 01920000 //;0017 ld	r9,r2		
      .INIT_02(256'h01920000_02940000_01930000_02b60000_07bb0200_01b60000_02a00000_04a00003),
// 07998300 //;0018 and	r9,r9,r8	
// b4f00012 //;0019 jz	cyc
// 02820000 //;001a st	r8,r2		
// 01950000 //;001b ld	r9,r5		
// 04a000ff //;001c ldl0	r10,0xff	
// 0799a400 //;001d xor	r9,r9,r10
// 02950000 //;001e st	r9,r5		
// b4f00012 //;001f jz	cyc
      .INIT_03(256'hb4f00012_02950000_0799a400_04a000ff_01950000_02820000_b4f00012_07998300),
// 01970000 //;0020 ld	r9,r7		
// 07990200 //;0021 inc	r9		
// 02970000 //;0022 st	r9,r7
// 04f00012 //;0023 jmp	cyc
      .INIT_04(256'h00000000_00000000_00000000_00000000_04f00012_02970000_07990200_01970000),
      .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .SRVAL(36'h000000000), .WRITE_MODE("WRITE_FIRST") ) RAM_L 
      (.ADDR(A[8:0]), 
                  .CLK(CLK), 
                  .DI(I[31:0]), 
                  .DIP({4'd0/*L, L, L, L*/}), 
                  .EN(CS), 
                  .SSR(1'b0/*L*/), 
                  .WE(WR), 
                  .DO(O[31:0]), 
                  .DOP());
   //GND  XLXI_7 (.G(L));
   //VCC  XLXI_9 (.P(H));
   //BUF  XLXI_10 (.I(CS), 
   //             .O(CSO));
endmodule