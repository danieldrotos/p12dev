module rfm2
  #(
    parameter WIDTH=32,
    parameter ADDR_SIZE=4
    )
   (
    input wire clk
    );
   
endmodule // rfm2
