module cpu2
  #(
    parameter WIDTH= 32,
    parameter ADDR_SIZE= 32
    )
  (
   // basic inputs
   input wire 		       clk,
   input wire 		       reset,
   // bus
   output wire [ADDR_SIZE-1:0] mbus_aout,
   input wire [WIDTH-1:0]      mbus_din,
   output wire [WIDTH-1:0]     mbus_dout,
   output wire 		       mbus_wen,
   // test
   input wire [3:0] 	       test_sel,
   output wire [WIDTH-1:0]     test_out,
   input wire [3:0] 	       test_rsel,
   output wire [WIDTH-1:0]     test_reg,
   output wire [2:0] 	       clk_stat
   );

   // internal signals
   wire [WIDTH-1:0] 	       ic;	// output of IC register
   wire [WIDTH-1:0] 	       pc;	// output of PC register 
   // phase signals
   wire 		       phf;	// fetch
   wire 		       phe;	// PC increment; execute
   wire 		       phm;	// memory r/w; link
   wire 		       phw;	// writeback
   // selected data as parameteres
   wire [WIDTH-1:0] 	       opa;
   wire [WIDTH-1:0] 	       opb;
   wire [WIDTH-1:0] 	       opd;
   // results
   wire [WIDTH-1:0] 	       res_alu;
   wire [7:0] 		       res_flags;
   wire [WIDTH-1:0] 	       res_call;
   wire [WIDTH-1:0] 	       res_ld;
   // selected data to use in writeback
   wire [3:0] 		       wb_address;
   wire [WIDTH-1:0] 	       wb_data;	// writeback data
   wire 		       wb_en;

   // scheduler generates phase signals
   schedm scheduler
     (
      .clk(clk),
      .reset(reset),
      .phf(phf),	// phase 1: FETCH (stores fetched code into IC reg)
      .phe(phe),	// phase 2: EXEC (signals go through ALU)
      .phm(phm),	// phase 3: MEM (LD/ST read/write)
      .phw(phw),	// phase 4: WRITEBACK (store back result to register)
      .clk_stat(clk_stat)
      );

   // FLAG register
   wire [7:0] 		       flags;
   wire 		       flag_c;
   wire 		       flag_s, flag_n;
   wire 		       flag_z;
   wire 		       flag_v, flag_o;
   wire 		       flag_p;
   wire 		       flag_u;
   wire 		       flag_wb_en;
   
   regm #(.WIDTH(8)) reg_flag
     (
      .clk(clk),
      .reset(reset/*1'b0*/),
      .cen(flag_wb_en),
      .din (res_flags),
      .dout(flags)
      );
   assign flag_c= flags[`CIDX];
   assign flag_s= flags[`SIDX];
   assign flag_z= flags[`ZIDX];
   assign flag_v= flags[`VIDX];
   assign flag_p= flags[`PIDX];
   assign flag_u= flags[`UIDX];
   assign flag_o= flag_v;
   assign flag_n= flag_s;
   assign flag_wb_en= ena & alu_wb_en & phw;

   // Instruction Register contains instruction code
   regm #(.WIDTH(WIDTH)) reg_ic
     (
      .clk(clk),
      .reset(reset),
      .cen(phf), // phe?
      .din(mbus_din),
      .dout(ic)
      );

   // pick parts of the IC
   wire 		       cond= ic[31:28];
   wire [2:0] 		       inst= ic[27:25];
   wire 		       inst_param= ic[24];
   wire [5:0] 		       alu_op= {ic[25:24],ic[19:16]};
   wire [3:0] 		       ra= ic[19:16];
   wire [3:0] 		       rb= ic[11:8];
   wire [3:0] 		       rd= ic[23:20];
   wire [15:0] 		       im16= ic[15:0];
   wire [23:0] 		       im24= ic[23:0];
   wire [19:0] 		       im20= ic[19:0];
   wire 		       u= ic[15];
   wire 		       p= ic[14];
   wire 		       w= ic[24];
   
   // decode instructions
   wire 		       inst_alu2= inst==0;
   wire 		       inst_alu1= inst==1;
   wire 		       inst_call= inst==2;
   wire 		       inst_ext = inst==3;
   wire 		       inst_st_r= inst==4;
   wire 		       inst_ld_r= inst==5;
   wire 		       inst_st_i= inst==6;
   wire 		       inst_ld_i= inst==7;
   wire 		       inst_alu;
   wire 		       inst_ld;
   wire 		       inst_st;
   wire 		       inst_mem;
   wire 		       inst_br;
   wire 		       inst_wb;
   assign inst_ld= inst_ld_r | inst_ld_i;
   assign inst_st= inst_st_r | inst_st_i;
   assign inst_mem= inst_st | inst_ld;
   assign inst_alu= inst_alu1 | inst_alu2;
   assign inst_br= inst_call | (inst_wb & (rd==4'd15));
   assign inst_wb= (inst_alu & alu_wb_en) |
		   inst_br |
		   inst_ld;

   // decode condition
   wire 		       ena;
   assign ena= (cond==4'h0)? 1 : // always
	       (cond==4'h1)? flag_z : // EQ
		     (cond==4'h2)? !flag_z : // NE
		     (cond==4'h3)? flag_c : // CS HS
		     (cond==4'h4)? !flag_c : // CC LO
		     (cond==4'h5)? flag_s : // MI
		     (cond==4'h6)? !flag_s : // PL
		     (cond==4'h7)? flag_o : // VS
		     (cond==4'h8)? !flag_o : // VC
		     (cond==4'h9)? flag_c & !flag_z : // HI
		     (cond==4'ha)? !flag_c | flag_z : // LS
		     (cond==4'hb)? !(flag_s ^ flag_o): // GE
		     (cond==4'hc)? flag_s ^ flag_o : // LT
		     (cond==4'hd)? !flag_z & !(flag_s ^ flag_o) : // GT
		     (cond==4'he)? flag_z | (flag_s ^ flag_o): // LE
		     (cond==4'hf)? 1 : // uncond
		     0;
   
   // ALU inst
   wire 		       alu_wb_en;
   wire 		       alu_flag_en;
   alu2 alu
     (
      // inputs
      .op(alu_op),
      .fi(flags),
      .bi(opb),
      .di(opd),
      .im(im16),
      // outputs
      .res(res_alu),
      .fo(res_flags),
      .wb_en(alu_wb_en),
      .flag_en(alu_flag_en)
      );

   // CALL inst
   wire [WIDTH-1:0] 	       aof_call_abs;
   wire [WIDTH-1:0] 	       aof_call_idx;
   wire [WIDTH-1:0] 	       sex_im20;
   wire 		       sof_im20= im20[19];
   assign sex_im20= {sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,sof_im20,im20};
   assign aof_call_abs= {8'b0, im24};
   assign aof_call_idx= opd+sex_im20;
   assign res_call= ic[24]?aof_call_idx:aof_call_abs;

   // Select data for write back
   assign wb_data= inst_alu?res_alu:
		   inst_call?res_call:
		   inst_ext?0:
		   inst_ld?mr_data:
		   inst_st?0:
		   0;
   assign wb_address= inst_call?4'd15:
		      rd;
   assign wb_en= ena & inst_wb & phw;

   // MEM inst (ld/st)
   wire [WIDTH-1:0] 	       mem_im_offset;
   assign mem_im_offset= {
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16[15],
			  im16
			  };
   wire [WIDTH-1:0] 	       aof_ldst;
   wire [WIDTH-1:0] 	       ldst_base;
   wire [WIDTH-1:0] 	       ldst_mod;
   wire [WIDTH-1:0] 	       opa_changed;
   wire [WIDTH-1:0] 	       ldst_offset;
   wire 		       up_down, pre_post;
   assign up_down= ic[26]?flag_u:u;
   assign pre_post= ic[26]?flag_p:p;
   assign ldst_mod= u?32'd1:32'hffffffff;
   assign opa_changed= opa+ldst_mod;
   assign ldst_base= pre_post?opa_changed:opa;
   assign ldst_offset= ic[26]?mem_im_offset:opb;
   assign aof_ldst= ldst_base+ldst_offset;

   // Register file
   rfm2 #(.WIDTH(WIDTH)) regs
     (
      .clk(clk),
      .reset(reset),
      .ra(ra),
      .rb(rb),
      .rd(rd),
      .rt(rt),
      .fn_inc_pc(phe),
      .fn_link(),
      .fn_ra_change(ena & inst_mem & w & phm),
      .fn_wb(ena & inst_wb & phw),
      .wb_data(wb_data),
      .ra_changed(opa_changed),
      .da(opa),
      .db(opb),
      .dd(opd),
      .dt(test_reg),
      .pc(pc)
      );
   
   // memory interface
   
   // handle input data lines
   wire 		       en_mr_data;
   assign en_mr_data= phm & inst_ld;
   // latched data read from memory
   reg [WIDTH-1:0] 	       mr_data;
   always @(posedge clk)
     begin
	if (en_mr_data)
	  mr_data<= mbus_din;
     end

   // produce address outputs
   wire [WIDTH-1:0] addr_phf;
   wire [WIDTH-1:0] addr_phe;
   wire [WIDTH-1:0] addr_phm;
   wire [WIDTH-1:0] addr_phw;

   assign addr_phf= pc;
   assign addr_phe= inst_ld?aof_ldst:pc;
   assign addr_phm= (inst_ld|inst_st)?aof_ldst:pc;
   assign addr_phw= (inst_br&ena)?wb_data:pc;
   assign mbus_aout= phf?addr_phf:
		     phe?addr_phe:
		     phm?addr_phm:
		     phw?addr_phw:
		     pc;

   // produce data outpouts   
   assign mbus_dout= opd;
   assign mbus_wen = ena & (phm/*|phe*/) & inst_st;

endmodule // cpu2
