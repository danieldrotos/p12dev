`timescale 1ns / 1ps

module mem(A, 
           CLK, 
           CS, 
           I, 
           WR, 
           CSO, 
           O);

    input [31:0] A;
    input CLK;
    input CS;
    input [31:0] I;
    input WR;
   output CSO;
   output [31:0] O;
   
   wire H;
   wire L;
   
   RAMB16_S36 #( 
      .INIT(36'h000000000), 
// //; SYMBOLS
// //; 0000c000 timer_ctrl
// //; 0000c001 timer_ar
// //; 0000c002 timer_cntr
// //; 0000c003 timer_stat
// //; 0000f000 display
// //; 0000f001 led
// //; 0000f002 portc
// //; 00000011 cyc
// //; CODE
// 00000000 //;0000 nop
// 0400c000 //;0001 ldl0	r0,timer_ctrl
// 0410c001 //;0002 ldl0	r1,timer_ar
// 0420c003 //;0003 ldl0	r2,timer_stat
// 0430c002 //;0004 ldl0	r3,timer_cntr
// 0440f000 //;0005 ldl0	r4,display
// 0450f001 //;0006 ldl0	r5,led
// 0460f002 //;0007 ldl0	r6,portc
      .INIT_00(256'h0460f002_0450f001_0440f000_0430c002_0420c003_0410c001_0400c000_00000000),
// 04700002 //;0008 ldl0	r7,2
// 04b00000 //;0009 ldl0	r11,0
// 04800000 //;000a ldl0	r8,0		
// 02850000 //;000b st	r8,r5
// 0590a120 //;000c ldl	r9,500000	
// 06900007 //;000d ldh	r9,500000
// 02910000 //;000e st	r9,r1
// 04a00003 //;000f ldl0	r10,3		
      .INIT_01(256'h04a00003_02910000_06900007_0590a120_02850000_04800000_04b00000_04700002),
// 02a00000 //;0010 st	r10,r0
// 07bb0200 //;0011 inc	r11		
// 02b60000 //;0012 st	r11,r6		
// 01830000 //;0013 ld	r8,r3		
// 02840000 //;0014 st	r8,r4		
// 01800000 //;0015 ld	r8,r0
// 04c0f003 //;0016 ldl0	r12,0xf003
// 028c0000 //;0017 st	r8,r12
      .INIT_02(256'h028c0000_04c0f003_01800000_02840000_01830000_02b60000_07bb0200_02a00000),
// 01820000 //;0018 ld	r8,r2		
// 07887300 //;0019 and	r8,r8,r7	
// b4f00011 //;001a jz	cyc
// 02720000 //;001b st	r7,r2		
// 01850000 //;001c ld	r8,r5		
// 049000ff //;001d ldl0	r9,0xff		
// 07889400 //;001e xor	r8,r8,r9
// 02850000 //;001f st	r8,r5		
      .INIT_03(256'h02850000_07889400_049000ff_01850000_02720000_b4f00011_07887300_01820000),
// 04f00011 //;0020 jmp	cyc
      .INIT_04(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_04f00011),
      .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000), 
      .SRVAL(36'h000000000), .WRITE_MODE("WRITE_FIRST") ) RAM_L 
      (.ADDR(A[8:0]), 
                  .CLK(CLK), 
                  .DI(I[31:0]), 
                  .DIP({4'd0/*L, L, L, L*/}), 
                  .EN(CS), 
                  .SSR(1'b0/*L*/), 
                  .WE(WR), 
                  .DO(O[31:0]), 
                  .DOP());
   //GND  XLXI_7 (.G(L));
   //VCC  XLXI_9 (.P(H));
   //BUF  XLXI_10 (.I(CS), 
   //             .O(CSO));
endmodule