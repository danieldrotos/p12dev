module rfm2
  #(
    parameter WIDTH=32
    )
   (
    input wire 	     clk,
    input wire 	     reset,
    input wire [3:0] ra,
    input wire [3:0] rb,
    input wire [3:0] rd,
    input wire [3:0] rt
    );
   
endmodule // rfm2
